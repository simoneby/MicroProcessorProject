module Datapath( // @[:@99.2]
  input   clock, // @[:@100.4]
  input   reset // @[:@101.4]
);
  initial begin end
endmodule

module Datapath( // @[:@238.2]
  input   clock, // @[:@239.4]
  input   reset // @[:@240.4]
);
  initial begin end
endmodule
